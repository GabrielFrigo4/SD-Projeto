package vending_machine is
    type state is (st0, st5, st10, st15, st20, st25, st30, st35, st40, st45, stcandy);
end package;

package body vending_machine is end package body;
