gabrielf@gabriel-vostro3520.1762:1754874173